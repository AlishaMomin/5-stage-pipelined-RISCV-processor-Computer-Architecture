module instruction_memory
(
    input [63:0] Inst_Address,
    output [31:0] Instruction
);
  reg [7:0] memory [131:0];
  initial begin  
//beq x11, x0, FinalExit
//100\\00000101\\1000110001100011
    memory[0] = 8'b01100011;
    memory[1] = 8'b10001100;
    memory[2] = 8'b00000101;
    memory[3] = 8'b00000100;  
    
//addi x4, x0, 0 
//imm|rs1|func3|rd|opcode
//000000000000|0000\\0|000|00100|0010011
    memory[4] = 8'b00010011;  
    memory[5] = 8'b00000010;
    memory[6] = 8'b00000000;
    memory[7] = 8'b00000000;

//beq x4, x11, Exit1
//10010110010\\00000110\\01100011
    memory[8] = 8'b01100011;
    memory[9] = 8'b00000110;
    memory[10] = 8'b10110010;
    memory[11] = 8'b00000100;   

//add x19, x0, x4
//0000000|00100|00000|000|10011|0110011
    memory[12] = 8'b10110011;
    memory[13] = 8'b00001001;
    memory[14] = 8'b01000000;
    memory[15] = 8'b00000000;
    
//beq x19, x11, Exit2
//10101110011000111001100011
    memory[16] = 8'b01100011;
    memory[17] = 8'b10001110;
    memory[18] = 8'b10111001;
    memory[19] = 8'b00000010; 

//slli x5, x4, 3
//000000000011|00100|001|00101|0010011  
    memory[20] = 8'b10010011;
    memory[21] = 8'b00010010;
    memory[22] = 8'b00110010;
    memory[23] = 8'b00000000;  
    
//slli x6, x19, 3 
//11|1001\\1|001|0011\\0|0010011
    memory[24] = 8'b00010011;
    memory[25] = 8'b10010011;
    memory[26] = 8'b00111001;
    memory[27] = 8'b00000000;  
   
//add x5, x5, x10 
//0000000|01010|00101|000|00101|0110011
    memory[28] = 8'b10110011;
    memory[29] = 8'b10000010;
    memory[30] = 8'b10100010;
    memory[31] = 8'b00000000; 
  
//add x6, x6, x10
//0000000|01010|00110|000|00110|0110011
    memory[32] = 8'b00110011;
    memory[33] = 8'b00000011;
    memory[34] = 8'b10100011;
    memory[35] = 8'b00000000;  
  
//ld x28, 0(x5)
//000000000000|00101|011|11100|0000011
    memory[36] = 8'b00000011;
    memory[37] = 8'b10111110;
    memory[38] = 8'b00000010;
    memory[39] = 8'b00000000;    
 
//ld x29, 0(x6)
//000000000000|00110|011|11101|0000011
    memory[40] = 8'b10000011;
    memory[41] = 8'b00111110;
    memory[42] = 8'b00000011;
    memory[43] = 8'b00000000; 
 
//bge x28, x29, iterate
//00000001110111100101110001100011
    memory[44] = 8'b01100011;
    memory[45] = 8'b01011100;
    memory[46] = 8'b11011110;
    memory[47] = 8'b00000001;    
    
//add x27, x0, x28
//        11100|00000|000|11011|0110011
//0000000|11100|00000|000|11011|0110011
    memory[48] = 8'b10110011;
    memory[49] = 8'b00001101;
    memory[50] = 8'b11000000;
    memory[51] = 8'b00000001;
    
//add x28, x0, x29
//func7|rs2|rs1|func3|rd|opcode
//0000000|11101|00000|000|11100|0110011
    memory[52] = 8'b00110011;
    memory[53] = 8'b00001110;
    memory[54] = 8'b11010000;
    memory[55] = 8'b00000001;   
 
//add x29, x0, x27
//0000000|1\\1011|0000\\0|000|11101|0110011
    memory[56] = 8'b10110011;
    memory[57] = 8'b00001110;
    memory[58] = 8'b10110000;
    memory[59] = 8'b00000001;    
  
//sd x28, 0(x5)
//00000|11100|00101|011|00000|0100011
    memory[60] =8'b00100011;
    memory[61] =8'b10110000;
    memory[62] =8'b11000010;
    memory[63] =8'b00000001;    
    
//sd x29, 0(x6)
//00000|11101|00110|011|00000|0100011
    memory[64] =8'b00100011;
    memory[65] =8'b00110000;
    memory[66] =8'b11010011;
    memory[67] =8'b00000001;    
    
//addi x19, x19, 1
//000000000001|10011|000|10011|0010011
    memory[68] =8'b10010011;
    memory[69] =8'b10001001;
    memory[70] =8'b00011001;
    memory[71] =8'b00000000;  
    
//beq x0, x0, Loop2
//11111100000000000000010011100011
    memory[72] =8'b11100011;
    memory[73] =8'b00000100;
    memory[74] =8'b00000000;
    memory[75] =8'b11111100;    
  
//addi x4, x4, 1
//imm|rs1|func3|rd|opcode
//000000000001|0010\\0|000|00100|0010011-------
    
    memory[76] =8'b00010011; 
    memory[77] =8'b00000010;
    memory[78] =8'b00010010;
    memory[79] =8'b00000000;
 
//beq x0, x0, Loop1
//00000000000000000000001011100011
    memory[80] =8'b11100011;
    memory[81] =8'b00001100;
    memory[82] =8'b00000000;
    memory[83] =8'b11111010;  
    
//beq x0, x0, FinalExit
//00000000000000000000001001100011
    memory[84] =8'b01100011;
    memory[85] =8'b00000010;  
    memory[86] =8'b00000000;
    memory[87] =8'b00000000; 
  
//FinalExit: nop
//00000000000000000000000000010011
    memory[88] =8'b00010011;
    memory[89] =8'b00000000;
    memory[90] =8'b00000000;
    memory[91] =8'b00000000;
  end
  assign Instruction = {memory[Inst_Address+3], memory[Inst_Address+2],
       memory[Inst_Address+1], memory[Inst_Address]}; 
endmodule